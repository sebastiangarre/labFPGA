library verilog;
use verilog.vl_types.all;
entity parte_e_vlg_vec_tst is
end parte_e_vlg_vec_tst;
