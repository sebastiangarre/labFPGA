library verilog;
use verilog.vl_types.all;
entity ejercicio2_vlg_vec_tst is
end ejercicio2_vlg_vec_tst;
