// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
// Created on Thu Nov 07 10:30:50 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module parte_e (
    reset,clock,sda,fin_dir,soy,fin_dato,
    hab_dir,hab_dato,ack);

    input reset;
    input clock;
    input sda;
    input fin_dir;
    input soy;
    input fin_dato;
    tri0 reset;
    tri0 sda;
    tri0 fin_dir;
    tri0 soy;
    tri0 fin_dato;
    output hab_dir;
    output hab_dato;
    output ack;
    reg hab_dir;
    reg hab_dato;
    reg ack;
    reg [5:0] fstate;
    reg [5:0] reg_fstate;
    parameter ocioso=0,start=1,guarda_dir=2,RorW=3,ackk=4,guarda_dato=5;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or sda or fin_dir or soy or fin_dato)
    begin
        if (reset) begin
            reg_fstate <= ocioso;
            hab_dir <= 1'b0;
            hab_dato <= 1'b0;
            ack <= 1'b0;
        end
        else begin
            hab_dir <= 1'b0;
            hab_dato <= 1'b0;
            ack <= 1'b0;
            case (fstate)
                ocioso: begin
                    if ((sda == 1'b0))
                        reg_fstate <= start;
                    else if ((sda == 1'b1))
                        reg_fstate <= ocioso;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= ocioso;

                    hab_dato <= 1'b0;

                    ack <= 1'b0;

                    hab_dir <= 1'b0;
                end
                start: begin
                    reg_fstate <= guarda_dir;

                    hab_dato <= 1'b0;

                    ack <= 1'b0;

                    hab_dir <= 1'b0;
                end
                guarda_dir: begin
                    if (((fin_dir == 1'b1) & (soy == 1'b0)))
                        reg_fstate <= ocioso;
                    else if ((fin_dir == 1'b0))
                        reg_fstate <= guarda_dir;
                    else if (((fin_dir == 1'b1) & (soy == 1'b1)))
                        reg_fstate <= RorW;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= guarda_dir;

                    hab_dato <= 1'b0;

                    ack <= 1'b0;

                    hab_dir <= 1'b1;
                end
                RorW: begin
                    reg_fstate <= ackk;

                    hab_dato <= 1'b0;

                    ack <= 1'b0;

                    hab_dir <= 1'b0;
                end
                ackk: begin
                    reg_fstate <= guarda_dato;

                    hab_dato <= 1'b0;

                    ack <= 1'b1;

                    hab_dir <= 1'b0;
                end
                guarda_dato: begin
                    if ((fin_dato == 1'b1))
                        reg_fstate <= ocioso;
                    else if ((fin_dato == 1'b0))
                        reg_fstate <= guarda_dato;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= guarda_dato;

                    hab_dato <= 1'b1;

                    ack <= 1'b0;

                    hab_dir <= 1'b0;
                end
                default: begin
                    hab_dir <= 1'bx;
                    hab_dato <= 1'bx;
                    ack <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // parte_e
