library verilog;
use verilog.vl_types.all;
entity ejercicio2_vlg_check_tst is
    port(
        output1         : in     vl_logic;
        output2         : in     vl_logic;
        output3         : in     vl_logic;
        output4         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ejercicio2_vlg_check_tst;
