-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Wed Nov 06 21:15:09 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Restador_Completo_4b IS 
	PORT
	(
		a0 :  IN  STD_LOGIC;
		b0 :  IN  STD_LOGIC;
		a1 :  IN  STD_LOGIC;
		b1 :  IN  STD_LOGIC;
		a2 :  IN  STD_LOGIC;
		b2 :  IN  STD_LOGIC;
		a3 :  IN  STD_LOGIC;
		b3 :  IN  STD_LOGIC;
		bin :  IN  STD_LOGIC;
		CLOCK :  IN  STD_LOGIC;
		bout :  OUT  STD_LOGIC;
		z3 :  OUT  STD_LOGIC;
		z2 :  OUT  STD_LOGIC;
		z1 :  OUT  STD_LOGIC;
		z0 :  OUT  STD_LOGIC
	);
END Restador_Completo_4b;

ARCHITECTURE bdf_type OF Restador_Completo_4b IS 

COMPONENT restador_completo
	PORT(in_a : IN STD_LOGIC;
		 in_b : IN STD_LOGIC;
		 in_bin : IN STD_LOGIC;
		 o_z : OUT STD_LOGIC;
		 o_bout : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	DFF_inst8 :  STD_LOGIC;
SIGNAL	DFF_inst9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	DFF_inst6 :  STD_LOGIC;
SIGNAL	DFF_inst11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	DFF_inst5 :  STD_LOGIC;
SIGNAL	DFF_inst12 :  STD_LOGIC;
SIGNAL	DFF_inst7 :  STD_LOGIC;
SIGNAL	DFF_inst10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_34 <= '1';
SYNTHESIZED_WIRE_35 <= '1';
SYNTHESIZED_WIRE_36 <= '1';
SYNTHESIZED_WIRE_37 <= '1';
SYNTHESIZED_WIRE_7 <= '1';
SYNTHESIZED_WIRE_10 <= '1';
SYNTHESIZED_WIRE_12 <= '1';
SYNTHESIZED_WIRE_38 <= '1';
SYNTHESIZED_WIRE_15 <= '1';
SYNTHESIZED_WIRE_16 <= '1';
SYNTHESIZED_WIRE_18 <= '1';
SYNTHESIZED_WIRE_39 <= '1';
SYNTHESIZED_WIRE_40 <= '1';
SYNTHESIZED_WIRE_41 <= '1';
SYNTHESIZED_WIRE_31 <= '1';
SYNTHESIZED_WIRE_33 <= '1';



b2v_inst : restador_completo
PORT MAP(in_a => DFF_inst8,
		 in_b => DFF_inst9,
		 in_bin => SYNTHESIZED_WIRE_0,
		 o_z => SYNTHESIZED_WIRE_14,
		 o_bout => SYNTHESIZED_WIRE_20);


PROCESS(CLOCK,SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
IF (SYNTHESIZED_WIRE_34 = '0') THEN
	DFF_inst10 <= '0';
ELSIF (SYNTHESIZED_WIRE_35 = '0') THEN
	DFF_inst10 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	DFF_inst10 <= b2;
END IF;
END PROCESS;


PROCESS(CLOCK,SYNTHESIZED_WIRE_35,SYNTHESIZED_WIRE_36)
BEGIN
IF (SYNTHESIZED_WIRE_35 = '0') THEN
	DFF_inst11 <= '0';
ELSIF (SYNTHESIZED_WIRE_36 = '0') THEN
	DFF_inst11 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	DFF_inst11 <= b1;
END IF;
END PROCESS;


PROCESS(CLOCK,SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
IF (SYNTHESIZED_WIRE_36 = '0') THEN
	DFF_inst12 <= '0';
ELSIF (SYNTHESIZED_WIRE_37 = '0') THEN
	DFF_inst12 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	DFF_inst12 <= b0;
END IF;
END PROCESS;


PROCESS(CLOCK,SYNTHESIZED_WIRE_7,SYNTHESIZED_WIRE_37)
BEGIN
IF (SYNTHESIZED_WIRE_7 = '0') THEN
	z0 <= '0';
ELSIF (SYNTHESIZED_WIRE_37 = '0') THEN
	z0 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	z0 <= SYNTHESIZED_WIRE_8;
END IF;
END PROCESS;


PROCESS(CLOCK,SYNTHESIZED_WIRE_10,SYNTHESIZED_WIRE_12)
BEGIN
IF (SYNTHESIZED_WIRE_10 = '0') THEN
	z1 <= '0';
ELSIF (SYNTHESIZED_WIRE_12 = '0') THEN
	z1 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	z1 <= SYNTHESIZED_WIRE_11;
END IF;
END PROCESS;


PROCESS(CLOCK,SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_15)
BEGIN
IF (SYNTHESIZED_WIRE_38 = '0') THEN
	z3 <= '0';
ELSIF (SYNTHESIZED_WIRE_15 = '0') THEN
	z3 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	z3 <= SYNTHESIZED_WIRE_14;
END IF;
END PROCESS;


PROCESS(CLOCK,SYNTHESIZED_WIRE_16,SYNTHESIZED_WIRE_18)
BEGIN
IF (SYNTHESIZED_WIRE_16 = '0') THEN
	z2 <= '0';
ELSIF (SYNTHESIZED_WIRE_18 = '0') THEN
	z2 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	z2 <= SYNTHESIZED_WIRE_17;
END IF;
END PROCESS;












PROCESS(CLOCK,SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_38)
BEGIN
IF (SYNTHESIZED_WIRE_38 = '0') THEN
	bout <= '0';
ELSIF (SYNTHESIZED_WIRE_38 = '0') THEN
	bout <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	bout <= SYNTHESIZED_WIRE_20;
END IF;
END PROCESS;








b2v_inst39 : restador_completo
PORT MAP(in_a => DFF_inst6,
		 in_b => DFF_inst11,
		 in_bin => SYNTHESIZED_WIRE_22,
		 o_z => SYNTHESIZED_WIRE_11,
		 o_bout => SYNTHESIZED_WIRE_23);


b2v_inst40 : restador_completo
PORT MAP(in_a => DFF_inst5,
		 in_b => DFF_inst12,
		 in_bin => bin,
		 o_z => SYNTHESIZED_WIRE_8,
		 o_bout => SYNTHESIZED_WIRE_22);


b2v_inst41 : restador_completo
PORT MAP(in_a => DFF_inst7,
		 in_b => DFF_inst10,
		 in_bin => SYNTHESIZED_WIRE_23,
		 o_z => SYNTHESIZED_WIRE_17,
		 o_bout => SYNTHESIZED_WIRE_0);


PROCESS(CLOCK,SYNTHESIZED_WIRE_39,SYNTHESIZED_WIRE_37)
BEGIN
IF (SYNTHESIZED_WIRE_39 = '0') THEN
	DFF_inst5 <= '0';
ELSIF (SYNTHESIZED_WIRE_37 = '0') THEN
	DFF_inst5 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	DFF_inst5 <= a0;
END IF;
END PROCESS;


PROCESS(CLOCK,SYNTHESIZED_WIRE_40,SYNTHESIZED_WIRE_39)
BEGIN
IF (SYNTHESIZED_WIRE_40 = '0') THEN
	DFF_inst6 <= '0';
ELSIF (SYNTHESIZED_WIRE_39 = '0') THEN
	DFF_inst6 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	DFF_inst6 <= a1;
END IF;
END PROCESS;


PROCESS(CLOCK,SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_40)
BEGIN
IF (SYNTHESIZED_WIRE_34 = '0') THEN
	DFF_inst7 <= '0';
ELSIF (SYNTHESIZED_WIRE_40 = '0') THEN
	DFF_inst7 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	DFF_inst7 <= a2;
END IF;
END PROCESS;


PROCESS(CLOCK,SYNTHESIZED_WIRE_41,SYNTHESIZED_WIRE_31)
BEGIN
IF (SYNTHESIZED_WIRE_41 = '0') THEN
	DFF_inst8 <= '0';
ELSIF (SYNTHESIZED_WIRE_31 = '0') THEN
	DFF_inst8 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	DFF_inst8 <= a3;
END IF;
END PROCESS;


PROCESS(CLOCK,SYNTHESIZED_WIRE_41,SYNTHESIZED_WIRE_33)
BEGIN
IF (SYNTHESIZED_WIRE_41 = '0') THEN
	DFF_inst9 <= '0';
ELSIF (SYNTHESIZED_WIRE_33 = '0') THEN
	DFF_inst9 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	DFF_inst9 <= b3;
END IF;
END PROCESS;


END bdf_type;