library verilog;
use verilog.vl_types.all;
entity Restador_Completo_vlg_vec_tst is
end Restador_Completo_vlg_vec_tst;
