library verilog;
use verilog.vl_types.all;
entity FPGAparteA_vlg_vec_tst is
end FPGAparteA_vlg_vec_tst;
