library verilog;
use verilog.vl_types.all;
entity Restador_Completo_vlg_check_tst is
    port(
        o_bout          : in     vl_logic;
        o_z             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Restador_Completo_vlg_check_tst;
