library verilog;
use verilog.vl_types.all;
entity Restador_Completo_4b_vlg_check_tst is
    port(
        bout            : in     vl_logic;
        z0              : in     vl_logic;
        z1              : in     vl_logic;
        z2              : in     vl_logic;
        z3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Restador_Completo_4b_vlg_check_tst;
