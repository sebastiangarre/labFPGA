library verilog;
use verilog.vl_types.all;
entity divisor_vlg_vec_tst is
end divisor_vlg_vec_tst;
