-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Thu Nov 07 10:31:47 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY parte_e IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        sda : IN STD_LOGIC := '0';
        fin_dir : IN STD_LOGIC := '0';
        soy : IN STD_LOGIC := '0';
        fin_dato : IN STD_LOGIC := '0';
        hab_dir : OUT STD_LOGIC;
        hab_dato : OUT STD_LOGIC;
        ack : OUT STD_LOGIC
    );
END parte_e;

ARCHITECTURE BEHAVIOR OF parte_e IS
    TYPE type_fstate IS (ocioso,start,guarda_dir,RorW,ackk,guarda_dato);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,sda,fin_dir,soy,fin_dato)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= ocioso;
            hab_dir <= '0';
            hab_dato <= '0';
            ack <= '0';
        ELSE
            hab_dir <= '0';
            hab_dato <= '0';
            ack <= '0';
            CASE fstate IS
                WHEN ocioso =>
                    IF ((sda = '0')) THEN
                        reg_fstate <= start;
                    ELSIF ((sda = '1')) THEN
                        reg_fstate <= ocioso;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ocioso;
                    END IF;

                    hab_dato <= '0';

                    ack <= '0';

                    hab_dir <= '0';
                WHEN start =>
                    reg_fstate <= guarda_dir;

                    hab_dato <= '0';

                    ack <= '0';

                    hab_dir <= '0';
                WHEN guarda_dir =>
                    IF (((fin_dir = '1') AND (soy = '0'))) THEN
                        reg_fstate <= ocioso;
                    ELSIF ((fin_dir = '0')) THEN
                        reg_fstate <= guarda_dir;
                    ELSIF (((fin_dir = '1') AND (soy = '1'))) THEN
                        reg_fstate <= RorW;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= guarda_dir;
                    END IF;

                    hab_dato <= '0';

                    ack <= '0';

                    hab_dir <= '1';
                WHEN RorW =>
                    reg_fstate <= ackk;

                    hab_dato <= '0';

                    ack <= '0';

                    hab_dir <= '0';
                WHEN ackk =>
                    reg_fstate <= guarda_dato;

                    hab_dato <= '0';

                    ack <= '1';

                    hab_dir <= '0';
                WHEN guarda_dato =>
                    IF ((fin_dato = '1')) THEN
                        reg_fstate <= ocioso;
                    ELSIF ((fin_dato = '0')) THEN
                        reg_fstate <= guarda_dato;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= guarda_dato;
                    END IF;

                    hab_dato <= '1';

                    ack <= '0';

                    hab_dir <= '0';
                WHEN OTHERS => 
                    hab_dir <= 'X';
                    hab_dato <= 'X';
                    ack <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
